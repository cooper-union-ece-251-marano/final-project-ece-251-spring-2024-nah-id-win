// //////////////////////////////////////////////////////////////////////////////////
// // The Cooper Union
// // ECE 251 Spring 2024
// // Engineer: Evan Rosenfeld, James Ryan
// // 
// //     Create Date: 2023-02-07
// //     Module Name: aludec
// //     Description: 32-bit RISC ALU decoder
// //
// // Revision: 1.0
// //
// //////////////////////////////////////////////////////////////////////////////////
// `ifndef ALUDEC
// `define ALUDEC

// `timescale 1ns/100ps

// module aludec
//     #(parameter n = 32)(
//     //
//     // ---------------- PORT DEFINITIONS ----------------
//     //

//     //
//     // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
//     //

// endmodule

// `endif // ALUDEC
