//////////////////////////////////////////////////////////////////////////////////
// The Cooper Union
// ECE 251 Spring 2024
// Engineer: Evan Rosenfeld, James Ryan
//
//     Create Date: 2024-05-02
//     Definitions file
//
// Revision: 1.0
//
//////////////////////////////////////////////////////////////////////////////////
`ifndef DEFINITIONS
`define DEFINITIONS

`define PC_REG 0
`define SP_REG 1
`define RA_REG 2
`define IM_REG 3
`define A_REG 4
`define X_REG 5
`define HI_REG 6
`define LO_REG 7
`define WORDSIZE 16
`define CW 4


`endif //DEFINITIONS
